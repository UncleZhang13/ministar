`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Myminieye
// Engineer: Nill
// 
// Create Date:   
// Design Name:  
// Module Name:  compare
// Project Name: 
// Target Devices: Gowin
// Tool Versions: 
// Description: 
//      
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

`define UD #1
module compare(
    input        clk,
    input [3:0]  sw,
    input [3:0]  ctrl,
    input        enter_trig,
    
    output       com_result
);

//==============================================================================
    //���浱ǰ���������룻
    reg [3:0] ctrl_1d;
    always @(posedge clk)
    begin
        if(enter_trig)
            ctrl_1d <= `UD ctrl;
    end

    assign com_result = (ctrl_1d == sw);
    
endmodule
